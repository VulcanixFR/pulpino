
module boot_code
(
		input  logic        CLK,
		input  logic        RSTN,

		input  logic        CSN,
		input  logic [9:0]  A,
		output logic [31:0] Q
	);

	const logic [0:547] [31:0] mem = {
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h00000013,
		32'h0100006F,
		32'h0100006F,
		32'h0080006F,
		32'h0040006F,
		32'h0000006F,
		32'h00000093,
		32'h00008113,
		32'h00008193,
		32'h00008213,
		32'h00008293,
		32'h00008313,
		32'h00008393,
		32'h00008413,
		32'h00008493,
		32'h00008513,
		32'h00008593,
		32'h00008613,
		32'h00008693,
		32'h00008713,
		32'h00008793,
		32'h00008813,
		32'h00008893,
		32'h00008913,
		32'h00008993,
		32'h00008A13,
		32'h00008A93,
		32'h00008B13,
		32'h00008B93,
		32'h00008C13,
		32'h00008C93,
		32'h00008D13,
		32'h00008D93,
		32'h00008E13,
		32'h00008E93,
		32'h00008F13,
		32'h00008F93,
		32'h00100117,
		32'hEF410113,
		32'h00000D17,
		32'h6DCD0D13,
		32'h00000D97,
		32'h6D4D8D93,
		32'h01BD5863,
		32'h000D2023,
		32'h004D0D13,
		32'hFFADDCE3,
		32'h00000513,
		32'h00000593,
		32'h074000EF,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h46811101,
		32'h45A14601,
		32'h09F00513,
		32'h00EFCE06,
		32'h051338A0,
		32'h00EF0400,
		32'h45813DE0,
		32'h00EF4501,
		32'h45813BE0,
		32'h00EF4501,
		32'h00284060,
		32'h04000593,
		32'h448000EF,
		32'h071347A2,
		32'hD5132190,
		32'h87A10187,
		32'hD7B3157D,
		32'h35331007,
		32'h886300A0,
		32'h670900E7,
		32'h8F990761,
		32'h00F037B3,
		32'h40F2953E,
		32'h80826105,
		32'h4505715D,
		32'hC4A2C686,
		32'hC0CAC2A6,
		32'hDC52DE4E,
		32'hD85ADA56,
		32'hD462D65E,
		32'hD06AD266,
		32'h268000EF,
		32'h45014585,
		32'h470000EF,
		32'h87936785,
		32'hC0FBBB87,
		32'h00010037,
		32'h47110001,
		32'h1A1027B7,
		32'hF0EFC3D8,
		32'hC911F63F,
		32'h00008537,
		32'h02400593,
		32'h74850513,
		32'h4A4000EF,
		32'h8537A001,
		32'h45C50000,
		32'h77050513,
		32'h494000EF,
		32'h46014681,
		32'h451945A1,
		32'h2CC000EF,
		32'h00EF4501,
		32'h64C13220,
		32'h45054581,
		32'h350000EF,
		32'h440514FD,
		32'h378000EF,
		32'h1DE38D65,
		32'h0637FE85,
		32'h06938000,
		32'h06130200,
		32'h45A13486,
		32'h07100513,
		32'h298000EF,
		32'h00EF4501,
		32'h64C12EE0,
		32'h85224581,
		32'h31C000EF,
		32'h00EF14FD,
		32'h8D653460,
		32'hFE851DE3,
		32'h45214581,
		32'h2B8000EF,
		32'h02000693,
		32'h45A14601,
		32'h0EB00513,
		32'h264000EF,
		32'h10000513,
		32'h2B8000EF,
		32'h45094581,
		32'h2E8000EF,
		32'h10000593,
		32'h00EF850A,
		32'h853732A0,
		32'h4CB20000,
		32'h051345D5,
		32'h44027845,
		32'h49C24C12,
		32'h4B724AD2,
		32'h3EC000EF,
		32'h45214581,
		32'h26C000EF,
		32'h07905F63,
		32'h642184A2,
		32'h0C334901,
		32'h8BB7409C,
		32'h04130000,
		32'h8A377E04,
		32'h6D050000,
		32'h00849613,
		32'h02000693,
		32'h051345A1,
		32'h00EF0EB0,
		32'h65211FA0,
		32'h250000EF,
		32'h45094581,
		32'h280000EF,
		32'h009C0533,
		32'h00EF65A1,
		32'h45992C20,
		32'h79CB8513,
		32'h394000EF,
		32'h00495513,
		32'h95224585,
		32'h388000EF,
		32'h00F97513,
		32'h95224585,
		32'h37C000EF,
		32'h45990905,
		32'h7A4A0513,
		32'h370000EF,
		32'h00EF94EA,
		32'h91E33AE0,
		32'h6441FB2C,
		32'h4485147D,
		32'h264000EF,
		32'h1DE38D61,
		32'h8537FE95,
		32'h45B50000,
		32'h7AC50513,
		32'h348000EF,
		32'h388000EF,
		32'h45214581,
		32'h1C4000EF,
		32'h07605F63,
		32'h84CE6421,
		32'h89B34901,
		32'h8BB7413A,
		32'h04130000,
		32'h8A377E04,
		32'h6A850000,
		32'h00849613,
		32'h02000693,
		32'h051345A1,
		32'h00EF0EB0,
		32'h65211520,
		32'h1A8000EF,
		32'h45094581,
		32'h1D8000EF,
		32'h00998533,
		32'h00EF65A1,
		32'h459921A0,
		32'h79CB8513,
		32'h2EC000EF,
		32'h00495513,
		32'h95224585,
		32'h2E0000EF,
		32'h00F97513,
		32'h95224585,
		32'h2D4000EF,
		32'h45990905,
		32'h7A4A0513,
		32'h2C8000EF,
		32'h00EF94D6,
		32'h11E33060,
		32'h8537FB2B,
		32'h05930000,
		32'h05130220,
		32'h00EF7BC5,
		32'h00EF2AE0,
		32'h77B72EE0,
		32'hA4231A10,
		32'h07930007,
		32'h80670800,
		32'h00010007,
		32'h00010001,
		32'h450140B6,
		32'h44964426,
		32'h59F24906,
		32'h5AD25A62,
		32'h5BB25B42,
		32'h5C925C22,
		32'h61615D02,
		32'h00008082,
		32'hFF010113,
		32'h00812423,
		32'h00000593,
		32'h00050413,
		32'h00F00513,
		32'h00112623,
		32'h00912223,
		32'h2B0000EF,
		32'h00000593,
		32'h00E00513,
		32'h2A4000EF,
		32'h00000593,
		32'h00D00513,
		32'h298000EF,
		32'h00000593,
		32'h00C00513,
		32'h28C000EF,
		32'h04805E63,
		32'h00100493,
		32'h00000593,
		32'h01000513,
		32'h278000EF,
		32'h04940463,
		32'h00000593,
		32'h00B00513,
		32'h268000EF,
		32'h00200793,
		32'h02F40A63,
		32'h00000593,
		32'h00000513,
		32'h254000EF,
		32'h00300793,
		32'h02F40063,
		32'h00048513,
		32'h00C12083,
		32'h00812403,
		32'h00412483,
		32'h00000593,
		32'h01010113,
		32'h2300006F,
		32'h00C12083,
		32'h00812403,
		32'h00412483,
		32'h01010113,
		32'h00008067,
		32'h00004837,
		32'hF0080813,
		32'h00869693,
		32'h02000713,
		32'h1A1027B7,
		32'h40B70733,
		32'h0106F6B3,
		32'h03F5F593,
		32'h00E51533,
		32'h00878813,
		32'h00C78713,
		32'h00B6E5B3,
		32'h01078793,
		32'h00A82023,
		32'h00C72023,
		32'h00B7A023,
		32'h00008067,
		32'h01059593,
		32'h10055533,
		32'h00A5E5B3,
		32'h1A1027B7,
		32'h00B7AA23,
		32'h00008067,
		32'h1A102737,
		32'h01070713,
		32'h00072783,
		32'hFF010113,
		32'h00F12623,
		32'h00C12783,
		32'h01051513,
		32'h1007D7B3,
		32'h00F56533,
		32'h00A12623,
		32'h00C12783,
		32'h01010113,
		32'h00F72023,
		32'h00008067,
		32'h00100793,
		32'h00858593,
		32'h00B795B3,
		32'h00A79533,
		32'h000017B7,
		32'hF0078793,
		32'h00F5F5B3,
		32'h0FF57513,
		32'h00A5E533,
		32'h1A1027B7,
		32'h00A7A023,
		32'h00008067,
		32'h1A1027B7,
		32'h0007A783,
		32'hFF010113,
		32'h00F12623,
		32'h00C12503,
		32'h01010113,
		32'h00008067,
		32'h4055D793,
		32'hFF010113,
		32'h7FF7F793,
		32'h01F5F593,
		32'h00F12423,
		32'h00058863,
		32'h00812783,
		32'h00178793,
		32'h00F12423,
		32'h00012623,
		32'h00C12683,
		32'h00812783,
		32'h1A102737,
		32'h02070813,
		32'h02F6DE63,
		32'h00072783,
		32'h4107D793,
		32'h0FF7F793,
		32'hFE078AE3,
		32'h00C12783,
		32'h00082583,
		32'h00C12683,
		32'h00279793,
		32'h00168693,
		32'h00D12623,
		32'h00C12603,
		32'h00812683,
		32'h1EB56023,
		32'hFCD646E3,
		32'h01010113,
		32'h00008067,
		32'h1A107737,
		32'h00470713,
		32'h00072603,
		32'h1A1007B7,
		32'h00266613,
		32'h00C72023,
		32'h00C78513,
		32'h08300713,
		32'h00E52023,
		32'h00478693,
		32'h0085D813,
		32'h00800713,
		32'h0FF5F593,
		32'h0106A023,
		32'h1CB7E02B,
		32'h0A700713,
		32'h00E7A023,
		32'h00300793,
		32'h00F52023,
		32'h0006A783,
		32'h0F07F793,
		32'h0027E793,
		32'h00F6A023,
		32'h00008067,
		32'h1A100737,
		32'h01470713,
		32'h02058863,
		32'h04000693,
		32'h00072783,
		32'h0207F793,
		32'hFE078CE3,
		32'h0015460B,
		32'h1A1007B7,
		32'hFFF58593,
		32'h00C7A023,
		32'hFFF68693,
		32'h00069663,
		32'hFC059CE3,
		32'h00008067,
		32'hFC059AE3,
		32'h00008067,
		32'h1A100737,
		32'h01470713,
		32'h00072783,
		32'h0407F793,
		32'hFE078CE3,
		32'h00008067,
		32'h1A1076B7,
		32'h0006A783,
		32'hFF010113,
		32'h00F12623,
		32'h00100793,
		32'h00C12703,
		32'h00A797B3,
		32'hFFF7C793,
		32'h00E7F7B3,
		32'h00F12623,
		32'h00C12783,
		32'h00A595B3,
		32'h00F5E533,
		32'h00A12623,
		32'h00C12783,
		32'h01010113,
		32'h00F6A023,
		32'h00008067,
		32'h4F525245,
		32'h53203A52,
		32'h736E6170,
		32'h206E6F69,
		32'h20495053,
		32'h73616C66,
		32'h6F6E2068,
		32'h6F662074,
		32'h0A646E75,
		32'h00000000,
		32'h64616F4C,
		32'h20676E69,
		32'h6D6F7266,
		32'h49505320,
		32'h0000000A,
		32'h79706F43,
		32'h20676E69,
		32'h74736E49,
		32'h74637572,
		32'h736E6F69,
		32'h0000000A,
		32'h636F6C42,
		32'h0000206B,
		32'h6E6F6420,
		32'h00000A65,
		32'h79706F43,
		32'h20676E69,
		32'h61746144,
		32'h0000000A,
		32'h656E6F44,
		32'h756A202C,
		32'h6E69706D,
		32'h6F742067,
		32'h736E4920,
		32'h63757274,
		32'h6E6F6974,
		32'h4D415220,
		32'h00000A2E,
		32'h33323130,
		32'h37363534,
		32'h42413938,
		32'h46454443,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000
	};

	logic [9:0] A_Q;

	always_ff @(posedge CLK)
	begin
		if (~RSTN)
			A_Q <= '0;
		else
			if (~CSN)
				A_Q <= A;
	end

	assign Q = mem[A_Q];

endmodule